library IEEE;
use ieee.std_logic_1164.all;

entity direccionar is

	port(
		numero_mezcladora: in std_logic_vector (1 downto 0);
		direccion: in std_logic_vector (7 downto 0);
		pertenece_grupo: in std_logic_vector (3 downto 0);
		M: out std_logic
	);

end entity;

architecture direction of direccionar is

component mux4a1_1bit is 
	port ( 
		control : in std_logic_vector (1 downto 0) ; 
		x0: in std_logic;
		x1: in std_logic;
		x2: in std_logic;
		x3: in std_logic;
		y:out std_logic
	); 
end component; 

signal p1, p2, p3, p4, M1, M2, M3, M4: std_logic;

begin

p1 <= (pertenece_grupo(0) and (not(direccion(2)) and not(direccion(3)))); --pertenece y envio a grupo1

p2 <= (pertenece_grupo(1) and (direccion(2) and not(direccion(3)))); --pertenece y envio a grupo2

p3 <= (pertenece_grupo(2) and (not(direccion(2)) and direccion(3))); --pertenece y envio a grupo3

p4 <= (pertenece_grupo(3) and (direccion(2) and direccion(3))); --pertenece y envio a grupo4

M1 <= (not(numero_mezcladora(0)) and not(numero_mezcladora(1)) and direccion(6) and not(direccion(0)) and not(direccion(1))) or direccion(5) or (direccion(4) and (p1 or p2 or p3 or p4));

M2 <= (numero_mezcladora(0) and not (numero_mezcladora(1)) and direccion(0) and not(direccion(1))) or direccion(5) or (direccion(4) and (p1 or p2 or p3 or p4));

M3 <= (not(numero_mezcladora(0)) and numero_mezcladora(1) and not(direccion(0)) and direccion(1)) or direccion(5) or (direccion(4) and (p1 or p2 or p3 or p4));

M4 <= (numero_mezcladora(0) and numero_mezcladora(1) and direccion(0) and direccion(1)) or direccion(5) or (direccion(4) and (p1 or p2 or p3 or p4));

MUXA: mux4a1_1bit
	port map( 
		control => numero_mezcladora, 
		x0 => M1,
		x1 => M2,
		x2 => M3,
		x3 => M4,
		y =>M
	); 


end architecture;